module myor(x, a, b);
output x;
input a, b;

or a0(x, a, b);
endmodule
