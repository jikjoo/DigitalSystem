module myxor(x, a, b);
output x;
input a, b;

xor a0(x, a, b);
endmodule