module mynand(x, a, b);
output x;
input a, b;

nand a0(x, a, b);
endmodule
