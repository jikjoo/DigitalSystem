module mynor(x, a, b);
output x;
input a, b;

nor a0(x, a, b);
endmodule