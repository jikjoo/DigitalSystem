module myand(x, a, b);
output x;
input a, b;

and a0(x, a, b);
endmodule
